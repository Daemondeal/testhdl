module Test;
initial begin
    $display("This is a test");
    $finish();
end
endmodule : Test

entity Test is
end Test;

architecture t of Test is
begin
  process
  begin
    report "Hello World";
    wait;
  end process;

end t;
